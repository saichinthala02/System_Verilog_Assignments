//--> Declaration of Ethernet packet.

class eth_pkt;
	static int count;
	rand bit[47:0]da;
	rand bit[15:0]len;
	rand byte payload[$];
		 bit[55:0]crc;

	function void print();
	//	count++;
		$display("-------------------");
	//	$display("Count:- %0d",count);
		$display("da=%0d",da);
		$display("len=%0d",len);
		$display("crc=%0d",crc);
		$display("payload=%p",payload);
	endfunction

	constraint len_c{
		len inside {[42:1500]};
		payload.size()==len;
	}
endclass

module top;
	eth_pkt pkt;
	initial begin
		pkt = new();
		repeat(10)begin
			pkt.randomize();
			pkt.count++;
			pkt.print();
		end
		$display("Total eth_pkt are %0d",pkt.count);
	end
endmodule

/* Output:-
# -------------------
# da=197270863703325
# len=753
# crc=0
# payload='{-51, -99, -18, -71, -68, -58, 20, 120, 111, 37, 31, -124, -1, 6, 115, 84, -91, 42, 118, 91, -108, 61, 19, 79, 111, -59, -30, 53, -61, -62, -40, 94, 109, -69, -94, 85, 35, -57, -70, -25, 121, -22, -38, -94, 81, -69, 98, 48, -57, -37, 123, 45, -55, -8, -91, -18, -79, 12, 72, -67, 66, -17, -124, -86, -38, 127, -35, -118, -48, 1, 102, 25, -55, 41, -82, 98, -6, -11, -29, 62, 44, 59, -94, -95, 50, -7, -76, -32, 7, 123, 22, -95, 26, -53, 16, 102, -69, -1, 104, -23, 80, -105, 81, -127, -31, 0, -47, -9, -79, -72, -88, -118, 63, -37, 69, 75, -102, -91, -40, 6, 104, 78, 90, -82, -66, 19, 110, 98, 57, 1, -94, -14, 15, 91, -107, -19, 109, -58, -97, -12, 107, -119, 105, -16, -6, -66, 27, 97, -52, 81, 124, 53, 8, 51, 38, -33, -52, -72, -101, -13, -29, 32, 77, -47, -86, -77, 78, 75, -121, -74, 7, -62, 54, -71, -60, -55, -72, -103, 50, 41, 0, 45, 79, 103, 115, -124, 98, 106, -1, -126, -87, -16, 25, -104, 46, 77, 126, -3, 60, -80, 77, -95, 106, -89, 58, -90, -92, 53, 27, -85, -55, -114, 9, 53, 21, -13, -22, -69, -128, -59, 90, -121, -47, 83, -67, 35, -41, -43, -108, 56, -84, 126, -79, -41, -119, -91, 95, 66, -31, -69, -99, -50, -119, 103, 13, 88, 82, -92, -11, -124, -46, 122, 68, 117, -63, 54, -7, 114, 78, -69, -120, 6, -78, -59, 87, 84, -40, -24, 122, 88, -106, -29, -37, 116, -60, -41, 28, -75, 98, -65, 47, -84, 78, -25, -5, -42, 18, -50, -5, 85, -106, 57, -104, -19, -91, 32, -39, 50, -36, 104, -62, 9, 105, -7, 101, 72, 66, -54, -13, -68, 60, -122, 27, 73, 81, 73, 50, 32, 95, -118, -76, 3, 118, -59, -101, -7, -124, 103, 40, 24, 107, -121, -110, 85, -4, 52, 113, 120, -4, -59, -56, 3, -12, 23, 7, 52, 34, -110, 41, 68, 36, 41, -20, 116, 67, 112, -8, 50, 20, -74, 7, -11, 15, -107, -44, 70, 118, 43, 71, -51, 43, 24, 32, 1, 119, 69, -31, 122, -74, 114, -59, 11, 25, 106, -122, -40, 58, -26, 76, -22, -50, -90, -75, 42, -125, -116, -28, -123, -70, -49, -55, -80, 127, -81, 30, 121, -6, -69, -72, -69, -116, 1, -11, 121, 23, 77, 5, -26, -114, 124, -49, -83, -95, -120, -110, -126, -4***trimmed
# -------------------
# da=58976385815933
# len=686
# crc=0
# payload='{85, 50, -88, 108, -47, -104, 104, -6, -90, 117, -49, -84, 47, 56, -114, 24, -102, 111, 15, -80, -28, 56, -54, 30, -128, -17, -3, 5, -63, -113, 39, -117, 113, -61, -22, 117, -70, -114, 46, 65, 69, -85, -32, -71, -125, 55, 81, -99, 91, -105, -110, -21, 111, -123, 110, -52, -85, 45, 81, -10, 87, 113, 101, -7, -66, -119, 33, 53, 50, -6, -73, -123, -120, -126, 23, 112, -42, 62, -70, -111, 59, 20, -96, 99, -127, 121, -41, -90, -62, -17, -121, 55, -31, -83, 105, 12, -35, 20, 65, 41, 85, -4, 125, 105, -84, 99, 100, -124, -71, 124, 40, -56, -122, -103, 77, 118, 16, -53, 96, -85, -101, -62, 76, 51, -98, -27, 29, -65, -109, -120, 96, -84, -56, 16, -103, -88, -44, -93, 107, -76, 98, 72, 70, 82, -42, -88, -23, 84, 40, 7, -39, 87, 40, -33, 55, -66, -57, 83, -125, 12, -20, -37, -55, -48, -43, -36, 81, 109, 110, -94, 114, 115, -34, 70, -110, -82, -59, -94, 2, 45, -42, -29, -91, -102, 125, -110, 102, -95, 121, 58, -65, -123, 60, -122, 88, -126, -25, 90, 82, 40, 26, -115, -40, -123, 2, -22, 61, 83, -69, 81, 121, -128, 33, -28, 112, -24, -114, 96, -30, -76, 47, 73, 32, -123, -85, -94, -7, 110, -19, 53, 112, -25, 83, 23, 97, 50, 87, -32, -75, -111, -103, 34, 36, -26, 25, 45, 48, -3, 121, -12, 12, 79, -65, -109, -27, -80, 15, 100, -31, -41, -45, 80, -47, -13, 103, -71, -126, 118, -115, -27, -44, -57, -25, -87, 98, 88, 74, -77, 22, -95, 78, 36, 46, 54, 28, -19, 74, 107, 14, 73, 123, 111, 92, -96, -52, 71, -114, -17, -39, 55, -113, 82, -34, 36, 32, 49, -5, 104, 95, 54, 88, -64, -61, -59, -65, 20, 6, 13, -12, -116, 34, -122, -85, -31, 53, -53, -97, -119, -70, 43, -117, 93, -111, 11, 109, 33, 22, 84, -103, -88, 66, 57, 49, 36, -61, -4, 125, -7, -69, 42, -35, -8, -93, -122, 63, -44, 60, -33, -45, -26, 55, 63, 98, -79, 31, 65, 91, 124, -36, 13, -63, 107, -99, 19, 110, -95, 98, -5, 57, -91, 50, -68, -6, -44, -51, 115, -23, 89, -24, -22, 58, 38, -106, -7, -56, -48, 35, -84, 64, -2, -12, 13, 15, -54, -117, -92, -110, 30, 118, 99, 22, 52, 47, 113, -77, -61, 90, 59, 121, 43, 30, -30, -***trimmed
# -------------------
# da=189399432218959
# len=1395
# crc=0
# payload='{60, 18, 68, -10, -14, -84, 42, 7, 71, 43, -117, 89, -80, -53, -60, 28, -54, -14, -33, -53, -15, -28, 29, -108, -31, -70, 87, -29, -45, 106, 118, 127, -111, -125, -2, 16, 118, -67, 65, 1, 63, 12, 53, -30, -8, 9, 83, 119, -85, -21, 15, -121, -96, 21, -26, -29, 30, 83, -16, 102, -30, -76, 108, -73, -65, 121, -117, -4, -46, 76, -59, -69, 107, 91, -102, -126, 83, -128, 104, -67, 49, 112, -96, 18, 17, -124, 119, 106, 78, -55, -48, 102, 64, 94, -117, 65, -53, 89, -98, -27, -126, 101, 45, 108, -8, -6, 121, 94, 42, -10, 110, 25, 99, -110, 113, -127, 123, -7, -44, -103, -112, -23, -89, 89, -17, 57, 26, 89, 29, -26, 122, -3, 5, 112, 2, 1, 39, 30, -107, -91, 121, 81, 98, 53, 11, -109, -8, -125, -60, 38, -21, 106, 71, -68, 56, -61, 82, -92, -2, 55, -80, 23, -35, 100, -36, 13, -66, -71, 7, -45, 115, -4, -61, -125, -80, -52, -71, 30, -85, -71, 97, 103, 98, -54, 15, 61, -56, -42, -22, -104, -42, -108, 117, -3, -75, -96, 1, 7, 114, -45, 53, -97, -17, 116, 104, -100, 34, 65, 32, -127, -57, 30, 111, -28, -112, 0, 119, 62, 12, 9, 77, 18, 42, 104, -1, -109, -44, -58, -26, -16, -83, -109, 118, -3, 16, 79, 99, -113, 68, 113, -35, 35, 8, 122, 87, 36, 74, 77, -17, 13, -117, -67, -58, 46, 111, 108, -18, -13, 124, 18, 84, -64, -117, -17, 40, -18, -92, -101, -126, -64, -36, -37, -6, -56, -90, -112, -104, 119, -2, 63, -39, 102, 49, -42, -72, -10, 10, -45, -21, 64, 85, -41, 30, 6, -14, -56, -72, 80, 59, 4, 29, -86, -8, 70, -106, 41, -123, 121, -119, 28, 29, 85, 57, 119, -3, -16, 23, -14, -95, -64, 61, -121, 71, 1, 90, -1, -120, 17, -51, 22, 76, 3, 51, -56, -69, 31, -65, -74, -10, 30, -12, 47, 120, -120, -126, -100, -49, -32, 29, 108, -17, -67, 121, -40, 52, 123, 96, 125, 49, 2, -9, -1, -80, -6, 45, -97, 122, -118, -30, -26, 13, -26, 113, -45, -63, -101, 77, -84, -79, -43, 101, -23, -126, -107, -34, -76, -72, -86, -63, 119, 71, 48, -69, 28, -59, 35, 84, -77, 13, -88, -20, -2, 66, -67, -69, -20, -93, -123, 122, -5, 96, 78, 123, -102, 92, -20, -57, 11, -68, 28, 117, 108, 19, -57, -11, -***trimmed
# -------------------
# da=27178819180587
# len=1249
# crc=0
# payload='{14, -112, -59, -38, -83, -20, -39, 68, 125, 97, 89, 37, 46, -35, -27, 24, -70, 2, 82, 15, -103, 10, -31, 59, 18, 109, -94, 13, -116, -84, -32, 81, -25, 24, 22, 9, -31, 41, 36, 19, -72, -111, 69, -14, -23, 43, -90, 64, -61, -75, -64, 111, -28, 103, -84, 102, -41, -104, 89, -108, -40, 119, 68, -64, -64, -75, 7, 84, 21, 43, -106, 63, -86, -34, -19, 76, 29, 72, 79, -39, -25, 57, 29, 100, 125, 88, -3, 41, -24, -111, 65, 22, 50, -45, -73, -127, -6, 38, 71, 19, 4, -33, 40, -94, 2, 7, 54, -13, 33, 59, -22, 127, 30, 27, -64, -40, -113, -107, 64, -63, 59, -23, -105, -108, -3, -7, 20, 10, 26, -111, -113, 59, 85, -16, 62, -13, -63, -118, -116, 34, 81, 49, 62, -44, -66, -111, 13, -14, 78, -103, -30, -11, 109, -109, 66, 73, 8, -29, -82, 72, -113, 43, -4, 7, 38, -40, -120, 45, -41, -70, -41, -76, 38, 2, -74, -127, -13, 83, -73, -46, 34, -92, -19, 89, 20, -91, -91, -47, -19, 25, -118, -105, -101, -37, 56, 105, 1, -35, -118, -39, -20, -118, -5, 81, -29, -126, -64, 67, 90, 32, -33, 127, 111, -3, 64, -11, 29, 28, 58, -58, 25, 25, -103, 102, 122, 36, -3, 5, 59, -87, -70, -39, -116, -118, 73, 85, 124, 53, 42, -105, 123, -91, 55, 98, 28, -15, 21, -112, -104, -6, 124, 63, 126, -35, -128, -84, 69, -45, -68, 99, 9, 29, 52, 79, 108, -35, 101, 95, -109, 27, 1, 123, -1, 99, 120, -87, -77, -63, 55, 40, 86, 74, -35, 84, 85, 7, -22, 101, 113, 21, -109, -21, 101, -46, -50, 45, -6, 94, -114, 62, -114, -126, -19, -62, 71, -43, -104, -31, 86, -73, 56, -66, 84, -58, 22, 127, -30, 55, -89, 71, -102, 89, 64, 87, 121, 122, 112, -9, -31, 45, 101, -77, 9, -56, 73, 116, -47, 43, -115, -125, 119, 28, 95, 17, 109, 17, -47, 95, -63, -28, 14, 50, -60, -1, -79, 34, 64, -46, 126, -73, 28, -67, -33, -53, 92, -82, 96, 81, 60, 12, -115, -73, 23, -62, 19, 51, 40, 50, -74, -29, -41, 11, -98, 69, -100, -78, -66, -10, -103, 31, 96, 58, 96, 8, 33, 45, 123, -115, 87, 72, -89, 15, 15, -46, -78, -70, 41, -71, 17, 5, 36, -81, 18, 25, 45, -95, 28, 117, 29, 124, 50, 102, -18, -23, 50, -82, 119, 118, -118, -110, -48***trimmed
# -------------------
# da=8372645406951
# len=594
# crc=0
# payload='{-57, 53, 5, 116, -103, -65, 33, 8, 105, 113, 13, 51, -1, 88, 17, -68, 63, -128, 19, 102, -1, 124, 97, 122, 103, 46, 16, 88, 79, -71, 118, 73, 107, -27, 17, -22, 42, -110, 67, 124, -44, 5, -98, 74, -28, -49, -73, -70, -54, -98, -78, -100, 84, -42, -119, 101, -3, -26, -27, -26, 66, -64, -99, 74, 76, 68, -22, 21, -71, -68, -1, -45, 102, 27, -125, 81, 30, 40, -82, 23, 6, -125, -20, -4, 112, 77, 11, 88, -106, 63, -106, -69, 90, -97, 74, 7, 38, -23, -64, 37, 6, 1, 59, -113, 16, 22, -67, 124, 121, -48, -74, 123, 118, -102, -18, 39, -14, -73, -32, 48, 69, -14, 41, 101, -32, -77, 43, -43, -25, -81, 23, -25, -67, 71, -41, -103, -22, -109, 59, 81, -104, 108, -24, 29, -33, -1, -105, 42, -63, -64, -31, -57, 35, 90, -114, 20, 49, 118, 43, 76, -6, 105, -110, 66, -123, 113, -56, -115, 126, -90, -1, -11, -12, 124, 88, -29, -52, 125, 71, 40, 97, -11, 79, -49, -97, 101, 111, -29, 88, 93, -123, -119, -82, 82, 103, 16, -55, 45, 42, 50, -13, -47, 97, 59, 44, -110, 76, -26, 111, 85, -56, -16, 97, -55, -39, -64, -84, 20, 127, 45, -89, 7, 108, -34, 41, 17, 33, -125, 123, 81, 41, -93, 106, 14, -128, 91, -83, -1, -70, 106, -28, 112, -82, -33, 112, 123, -75, -73, -91, 88, 125, -73, 22, 22, -114, 62, 95, -113, -86, -36, -53, -122, -108, -84, 92, 98, -99, -114, -127, -14, -106, -4, -18, 25, -34, 103, 115, 57, 104, -105, 44, 78, -79, -88, -51, -24, 117, 83, 81, -127, -69, 85, 76, 66, -109, 84, 127, 63, 100, 54, 101, -64, 69, -4, 70, -12, 44, -14, 30, -109, 32, -50, 74, 10, 102, -120, 45, 65, 112, -93, -32, -27, -78, 96, -104, 48, -72, 92, -74, 123, 109, 77, 117, -48, -42, -84, -94, -114, 33, 76, -89, -47, 19, 64, 105, -94, -69, -66, 76, -37, 108, -88, -90, 119, 60, -61, -57, 65, 116, -4, 18, -108, 68, 18, 97, -45, -34, 115, 14, 14, -72, 95, 27, -128, 100, -66, 44, 26, 57, -45, -70, 12, 86, -95, -103, 92, 27, -19, 101, -28, -82, 90, 26, -82, -5, -47, 4, 121, -74, -53, 51, 67, -123, -28, 17, 14, 1, 80, -64, 49, 102, 78, 0, 44, -51, -86, -105, 126, 45, 25, 92, -128, -119, -15, -112, -81,***trimmed
# -------------------
# da=106330588620994
# len=647
# crc=0
# payload='{28, 99, 105, -30, 81, 13, 94, -22, 125, 88, 127, 112, -117, -88, 28, -80, -76, 43, -22, 98, 75, -106, -125, -100, 56, 8, -92, 42, -21, 83, 38, -98, 31, -13, -96, -41, -53, 74, -111, -73, -31, 49, -100, -10, -10, 106, -6, 42, -106, -104, 32, 99, 74, -69, -128, -11, -117, 30, -45, 64, 16, -30, 88, -27, 32, 86, 64, 81, -80, -118, -121, -46, 75, 42, -108, 125, -47, -63, -57, 18, -99, 123, 107, 36, -56, -87, 47, 127, -106, -70, -43, 71, 18, 16, 84, 67, 55, -103, 55, -50, 99, 14, -46, 106, 78, -113, -5, 43, 21, 105, 78, -25, -63, 85, -82, -119, 71, 91, 20, -90, -9, 63, 109, -23, 72, -74, 111, -125, 92, 111, -67, -26, -112, 46, -104, -18, -117, 80, 9, 106, -118, 92, -39, -97, 113, -96, -114, 106, -37, -65, 30, 71, 96, -53, 35, 15, -33, -85, 69, -35, 11, -35, 3, -7, 30, -63, -105, -19, -102, -33, 38, 4, -58, 2, 46, 118, -30, -9, 27, -17, 23, 7, 14, 96, 113, 32, 121, 123, -81, -115, -17, 124, 119, -62, 97, -47, -3, 88, 43, -120, -44, -3, 46, 39, -54, 24, 51, 22, 103, 27, 95, -102, 114, 50, -59, 100, 29, 67, -21, -125, 78, 120, -101, 69, -3, -52, 115, -17, 4, 22, 100, 70, 16, -71, -6, 101, 107, -86, 76, -84, -26, 80, 62, -13, -52, -88, 1, 91, 63, -35, 5, 93, -68, -41, -52, -75, 72, -34, 117, 34, -37, -82, -30, -70, -120, 105, -42, 101, 124, -80, -18, 64, 27, -74, -56, 127, 83, -47, -20, -49, 4, 59, -91, -42, 55, -14, 12, 56, 127, 92, -82, 26, -98, -112, -63, 38, 44, 110, 113, -61, -55, 111, -113, 66, -117, -16, -104, -19, 121, 108, -99, -23, 99, -114, -41, -41, 127, -107, 46, -99, 80, -20, -22, 39, 86, -24, 89, -64, -12, 29, -25, -117, 108, -86, 18, 23, -59, -120, 69, -109, -97, 99, -81, 26, 79, 97, -116, 120, 5, 73, 22, -4, 50, -122, 96, 73, -117, -19, 90, 2, -26, -86, -15, 66, -107, -30, -74, 88, 54, 84, 32, 96, 54, 13, -40, -116, -92, 103, -54, -103, 49, 106, -59, -40, 56, 0, 122, 21, 0, -13, 108, 119, -28, -61, -121, 17, -12, -89, -4, 59, -19, 117, 41, 97, 25, 55, 33, 111, -103, -73, 1, 101, 125, -108, -5, 31, -104, 2, -128, -15, 75, -40, -121, -67, -12, -45, ***trimmed
# -------------------
# da=26738940385388
# len=1253
# crc=0
# payload='{-58, 75, -79, -102, -105, 28, 70, 52, 14, -100, -47, 79, -19, -109, -66, 41, -105, 25, 49, -56, -45, 78, 94, 60, -125, -101, 105, 91, 7, 83, 37, -39, -128, -68, 55, -52, -93, -119, 20, 97, 41, 44, 7, -71, 32, 82, 47, -33, -63, 95, 58, -19, 69, 87, -108, -92, -66, -76, -88, 27, -31, -30, 26, 113, 92, 33, 33, -86, 100, -31, -9, 78, 90, -114, 93, -81, 121, 30, 106, -66, -34, -38, 67, 101, 15, 89, -87, -72, 39, 88, -116, 71, -76, -89, -27, 62, -87, 15, 111, 103, -117, 119, -60, -21, 2, 35, 96, -91, -73, -38, -61, -101, -47, 79, 68, 8, -33, 10, -115, -17, 106, -111, -124, -72, -11, -102, -64, -92, 111, 106, -3, 67, 84, 6, -7, -10, 40, -50, 35, 21, -107, -31, -9, -26, 6, -101, -93, 64, -103, -72, -59, 99, 72, 65, 63, -114, 27, -46, -8, -61, -4, -101, 62, 125, 14, 21, 39, -18, -116, -80, -24, -92, 91, 9, 4, -26, -47, 4, -15, -65, -124, 70, 9, -48, 84, -82, -119, 49, -42, -85, -117, -103, -9, -115, -91, 55, 122, 61, 48, 38, 112, -36, -118, 125, 30, -87, -2, -118, -31, -72, -20, 43, 96, -69, 4, -78, -67, -100, 8, 42, -45, 39, -110, -6, 81, 60, 36, 116, -10, -83, -108, -120, -118, 112, -108, 67, 74, 38, -85, -44, 1, -79, -23, 78, -65, -73, -20, -54, -68, -85, 38, 9, -47, -103, 74, 87, 62, 39, 127, 69, -45, 7, -95, 85, -86, 118, 20, -58, -113, 110, -76, 100, 65, -123, 73, 27, -75, 36, 83, -20, -90, 118, 15, 72, -101, -58, 16, -37, -49, 77, -43, 102, -123, 70, 38, 24, -47, -63, 107, 89, -56, -107, -89, 28, 16, -111, 33, 9, -65, 91, -40, 32, -25, 69, 90, 11, 26, 117, 92, -61, 20, 73, 63, 3, -5, 108, -29, -112, 24, -12, -65, -86, -9, 75, -122, 61, 24, 78, -97, 23, 48, -65, 113, 46, 51, -49, -29, -114, -49, -10, 103, 1, -78, -31, -79, 90, 117, -87, 10, 110, 24, 105, 84, -56, -72, 82, -124, -115, 17, 45, 85, -111, 13, -39, -7, -76, 39, 12, -113, -5, 15, -31, 89, 91, 37, -50, 92, -71, -110, -104, 29, -25, -90, 94, -51, -40, -69, 38, -100, 82, 55, -69, -9, -68, 69, -13, -99, 61, -66, 73, -3, -78, -42, 56, -43, 53, -38, 108, 84, -126, 90, -76, 52, 53, 13, -60, 42, 94, 65, ***trimmed
# -------------------
# da=133456015071495
# len=756
# crc=0
# payload='{73, -120, 62, 34, -17, -78, 16, 93, -26, 24, -76, 118, 54, -85, -93, -60, -16, -89, 81, 55, 119, 43, 76, -89, 96, -115, 19, -105, 83, 113, 42, 100, 46, 24, -53, 16, -111, 52, -17, 126, 76, -45, 101, 63, 118, 83, -119, 104, -5, -3, 47, -127, 18, -13, 14, -10, 20, 90, -127, -61, -119, 11, 40, -108, 60, 92, 5, 84, -47, 48, 5, -48, -115, 125, 71, 110, 102, -11, -120, 32, -87, -91, -82, 10, -128, 20, -28, 0, -128, 70, 75, 114, 116, -1, 82, 52, 34, -101, -125, -62, 111, -77, 9, 127, -7, -10, -73, -63, 90, -31, 119, 49, -86, -63, -49, -26, 43, 108, -107, -4, -47, -73, 4, -105, 51, -123, 100, 87, 118, -16, 54, -10, -8, 69, -95, -34, 86, 127, 56, -54, -128, 18, -25, -114, 83, 29, -97, -110, 19, 20, -28, -109, 125, -89, 13, 32, 75, 47, 34, -42, -85, 24, 20, 96, -40, 97, -122, 15, 12, -56, 18, 120, -22, 56, -61, -46, -108, -36, 77, 93, 79, 8, 6, -19, -111, -87, -72, -58, -23, -55, -118, 87, -79, -85, -102, 107, -42, -2, 65, 64, -93, 8, 82, -95, -19, -51, -124, 86, 36, -72, 30, -10, 4, -51, -124, -36, 21, -87, 78, 15, -116, 70, 127, -105, -32, -94, 103, 28, -66, 3, -119, 38, -63, -10, 21, 91, -69, -98, -39, -73, 122, -15, -118, -76, -67, 109, -9, 86, -125, -6, 48, 75, 6, 81, -96, -99, 44, -38, -92, 100, -5, -118, 81, -56, -100, 89, -26, -72, 45, 61, 39, -18, -73, -89, -8, -20, 48, 125, -3, -127, -123, -116, 79, -63, 21, 43, -34, -106, -31, -109, -106, -88, 9, 64, 27, -65, -62, -43, -9, -8, -56, -74, 46, -56, -126, 35, 15, 61, -53, -88, 97, 48, 121, -74, 50, 121, -79, -50, 106, 111, 105, 58, 79, 70, 33, -48, 63, 36, -58, 23, 77, -70, -128, -102, -92, -22, -89, 0, 69, 106, -33, -98, 20, -125, -123, -55, -20, 115, 39, 80, -98, -29, -90, 51, -117, -65, 125, 59, 54, 69, 38, -103, 10, 5, 114, 91, 31, 14, 42, -94, -126, 53, -22, 25, 30, -49, 115, 110, 65, 125, 118, 6, -123, -48, 73, -35, -39, -70, 9, 106, 40, 114, 125, -89, -38, 36, 97, -66, -30, -81, 59, -65, 15, -74, 5, 46, -122, 0, 99, -107, 41, -119, -7, -27, 82, -11, 58, -31, -119, 48, -86, 103, 55, -80, 101, -46, 60,***trimmed
# -------------------
# da=181654478713871
# len=822
# crc=0
# payload='{-5, 104, -42, 77, -120, 32, -62, 57, -13, 93, -95, -59, 98, 124, -77, -40, 75, 84, 79, -109, 98, 52, 78, -45, -42, 109, 17, 5, -109, -37, 86, 53, -116, 39, 93, -44, 110, -42, 5, 66, -90, 3, -51, 78, 40, -21, 50, 71, -85, -2, -62, -79, -6, 105, -89, 119, -73, 111, -17, 55, 7, 60, -24, -83, -103, -22, -91, 65, -67, 12, 51, 75, -25, -14, -70, -51, -79, -59, -91, -11, 101, -70, 13, -115, -45, 49, -73, -42, -90, -56, 83, 85, 42, -33, 95, 60, -89, -110, -122, -126, -88, -81, -1, -65, 75, -7, 99, -88, 22, 101, -2, -69, 51, -7, -105, 12, 109, 49, -103, 0, 71, 113, 80, -107, 60, -120, -23, -91, 60, -74, -111, -60, -16, 89, 45, -94, 110, -60, -65, 55, -112, -60, -50, -82, 83, -51, -14, 82, -36, 58, -110, 59, 65, 74, -114, 120, -5, 80, -6, 86, -14, 37, -16, -14, 39, 55, -117, -92, -8, -83, 51, -111, 11, -82, 0, -115, 41, -46, -33, -93, 14, -3, 107, 31, 116, -70, -99, 103, 56, -45, 13, -61, -54, 45, -36, 43, 89, 116, 22, 47, 88, 34, 41, -75, -91, -126, 93, -43, 94, 7, -102, -116, 108, -53, -75, -81, 123, -28, -42, 44, -53, -118, 62, 25, 32, -116, 36, 42, -16, -114, -21, 106, 29, 76, 47, 91, -122, 6, -127, 5, 18, -25, -41, -57, 76, 77, 92, 9, -56, -112, -121, 17, 71, -109, -108, -88, 90, 83, -76, -91, 121, 110, -28, 17, -49, 119, 90, -96, 64, -27, -120, 52, 28, 68, 53, -37, -38, 68, 74, 65, -29, 57, -83, -41, -1, 16, -61, -68, -61, 93, -18, -110, -14, 80, 71, 123, -74, 22, 121, 42, -67, -123, -57, 96, 50, 28, -116, 67, -31, 0, 90, 15, -15, -40, 43, -89, -40, -17, 122, -17, -36, 21, 43, -73, 93, -8, -80, -33, -63, 111, 76, 70, 43, -53, 50, 27, 79, 19, -87, -2, 39, 97, 91, -71, -118, -8, -85, 120, 36, 28, -8, -100, -66, 9, 124, -62, 20, 82, 7, -119, 114, -35, 63, -87, -56, 13, 28, -116, 14, -2, -125, 36, 64, -85, 65, 12, 121, -115, -32, 34, 45, 44, 29, 38, 114, -2, 98, -44, 78, -10, -116, 58, 38, 16, -64, -86, -110, 15, 90, -110, 18, 84, -7, -100, 96, 42, 81, 116, 123, 68, 111, -2, -92, -86, -6, 76, -41, -37, -123, -123, 81, -124, -12, 39, 44, -93, 63, -13, -123, 30, 1***trimmed
# -------------------
# da=106442807273886
# len=81
# crc=0
# payload='{-4, 48, -121, 89, -4, -90, -124, -64, 110, -56, -57, 8, 49, -81, -95, 27, -33, 57, 97, -23, -77, -90, -24, 20, 45, -10, 34, -65, 9, 2, 90, 35, -47, -123, 37, -121, 74, -32, -123, -111, -118, 4, -85, -22, 116, -106, -48, -73, -47, -15, 24, -114, 25, -69, 124, -35, -119, 35, -107, -116, -102, 67, -82, -98, 48, 52, -121, -2, -81, -81, 24, 97, -76, -120, -11, -38, 58, 13, -52, -4, -34}
# Total eth_pkt are 10
*/
