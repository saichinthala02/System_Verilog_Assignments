//--> Q17. Operators.
module top;
	int a,c,b;
	initial begin
		a=10;
		b=12;
		$display("-----------------------------------------------");
		$display("--------> a=b <-------- ");
		$display("A:- %0d || B:- %0d",a,b);
		a=b;
		$display("A:- %0d || B:- %0d",a,b);
		$display("-----------------------------------------------");
		$display("--------> a+=b <-------- ");
		a=06;
		b=07;
		$display("A:- %0d || B:- %0d",a,b);
		a+=b;
		$display("A:- %0d || B:- %0d",a,b);
		$display("-----------------------------------------------");
		$display("--------> a-=b <-------- ");
		a=12;
		b=12;
		$display("A:- %0d || B:- %0d",a,b);
		a-=b;
		$display("A:- %0d || B:- %0d",a,b);
		$display("-----------------------------------------------");
		$display("--------> a*=b <-------- ");
		a=03;
		b=03;
		$display("A:- %0d || B:- %0d",a,b);
		a*=b;
		$display("A:- %0d || B:- %0d",a,b);
		$display("-----------------------------------------------");
		$display("--------> a/=b <-------- ");
		a=14;
		b=07;
		$display("A:- %0d || B:- %0d",a,b);
		a/=b;
		$display("A:- %0d || B:- %0d",a,b);
		$display("-----------------------------------------------");
		$display("--------> a%%=b <-------- ");
		a=12;
		b=4;
		$display("A:- %0d || B:- %0d",a,b);
		a%=b;
		$display("A:- %0d || B:- %0d",a,b);
		$display("-----------------------------------------------");
		$display("--------> a&=b <-------- ");
		a=10;
		b=12;
		$display("A:- %b || B:- %b",a,b);
		a&=b;
		$display("A:- %b || B:- %b",a,b);
		$display("-----------------------------------------------");
		$display("--------> a|=b <-------- ");
		a=10;
		b=12;
		$display("A:- %b || B:- %b",a,b);
		a|=b;
		$display("A:- %b || B:- %b",a,b);
		$display("-----------------------------------------------");
		$display("--------> a^=b <-------- ");
		
		a=10;
		b=12;

		$display("A:- %b || B:- %b",a,b);
		a^=b;
		$display("A:- %b || B:- %b",a,b);
		$display("-----------------------------------------------");
		$display("--------> a<<=2 <-------- ");

		a=7;
		$display("A:- %b",a);
		a<<=2;
		$display("A:- %b",a);
		$display("-----------------------------------------------");
		$display("--------> a>>=2 <-------- ");
		a=7;
		$display("A:- %b",a);
		a>>=2;
		$display("A:- %b",a);
		$display("-----------------------------------------------");
		$display("--------> a<<<=2 <-------- ");
		a=-07;
		$display("A:- %b",a);
		a<<<=2;
		$display("A:- %b",a);
		$display("-----------------------------------------------");
		$display("--------> a>>>=2 <-------- ");
		a=-07;
		$display("A:- %b",a);
		a>>>=2;
		$display("A:- %b",a);
		$display("-----------------------------------------------");
		a= 30; b=60;
		c= a+b;
		$display("\t--> ADD A:- %0d | B:- %0d || C:- %0d",a,b,c); 
		a= 60; b=20;
		c= a-b;
		$display("\t--> SUB A:- %0d | B:- %0d || C:- %0d",a,b,c); 
		a= 30; b=60;
		c= a*b;
		$display("\t--> MUL A:- %0d | B:- %0d || C:- %0d",a,b,c); 
		a= 30; b=05;
		c= a/b;
		$display("\t--> DIV A:- %0d | B:- %0d || C:- %0d",a,b,c); 
		a= 30; b=05;
		c= a%b;
		$display("\t--> MOD A:- %0d | B:- %0d || C:- %0d",a,b,c); 
		a= 2; b=12;
		c= a**b;
		$display("\t--> POW A:- %0d | B:- %0d || C:- %0d",a,b,c);
		$display("-----------------------------------------------");
		a= 4'b1011;
		b= 4'b0011;
		c= a&b;
		$display("\t--> AND A:- %0b B:- %0b C:- %0b",a,b,c); 
		c= a|b;
		$display("\t--> OR A:- %0b B:- %0b C:- %0b",a,b,c); 
		c= ~(a&b);
		$display("\t--> NAND A:- %0b B:- %0b C:- %0b",a,b,c); 
		c= ~(a|b);
		$display("\t--> NOR A:- %0b B:- %0b C:- %0b",a,b,c); 
		c= a^b;
		$display("\t--> XOR A:- %0b B:- %0b C:- %0b",a,b,c); 
		c= ~(a^b);
		$display("\t--> XNOR A:- %0b B:- %0b C:- %0b",a,b,c); 
		c = ~a;
		$display("\t--> NOT A:- %0b C:- %0b",a,c); 
		c = ~b; 
		$display("\t--> NOT B:- %0b C:- %0b",b,c);
		$display("-----------------------------------------------");
		a=4'b1000;
		b=4'b0000;
		c= a&&b;
		$display("\t--> LOGICAL_AND A:- %0b B:- %0b C:- %0b",a,b,c); 
		c= !(a&&b);
		$display("\t--> LOGICAL_!AND A:- %0b B:- %0b C:- %0b",a,b,c); 
		c= a||b;
		$display("\t--> LOGICAL_OR A:- %0b B:- %0b C:- %0b",a,b,c); 
		c= !(a||b);
		$display("\t--> LOGICAL_!OR A:- %0b B:- %0b C:- %0b",a,b,c);
		$display("-----------------------------------------------");
	end
endmodule

/* Output:-
# Start time: 19:53:10 on Nov 04,2025
# -----------------------------------------------
# --------> a=b <-------- 
# A:- 10 || B:- 12
# A:- 12 || B:- 12
# -----------------------------------------------
# --------> a+=b <-------- 
# A:- 6 || B:- 7
# A:- 13 || B:- 7
# -----------------------------------------------
# --------> a-=b <-------- 
# A:- 12 || B:- 12
# A:- 0 || B:- 12
# -----------------------------------------------
# --------> a*=b <-------- 
# A:- 3 || B:- 3
# A:- 9 || B:- 3
# -----------------------------------------------
# --------> a/=b <-------- 
# A:- 14 || B:- 7
# A:- 2 || B:- 7
# -----------------------------------------------
# --------> a%=b <-------- 
# A:- 12 || B:- 4
# A:- 0 || B:- 4
# -----------------------------------------------
# --------> a&=b <-------- 
# A:- 00000000000000000000000000001010 || B:- 00000000000000000000000000001100
# A:- 00000000000000000000000000001000 || B:- 00000000000000000000000000001100
# -----------------------------------------------
# --------> a|=b <-------- 
# A:- 00000000000000000000000000001010 || B:- 00000000000000000000000000001100
# A:- 00000000000000000000000000001110 || B:- 00000000000000000000000000001100
# -----------------------------------------------
# --------> a^=b <-------- 
# A:- 00000000000000000000000000001010 || B:- 00000000000000000000000000001100
# A:- 00000000000000000000000000000110 || B:- 00000000000000000000000000001100
# -----------------------------------------------
# --------> a<<=2 <-------- 
# A:- 00000000000000000000000000000111
# A:- 00000000000000000000000000011100
# -----------------------------------------------
# --------> a>>=2 <-------- 
# A:- 00000000000000000000000000000111
# A:- 00000000000000000000000000000001
# -----------------------------------------------
# --------> a<<<=2 <-------- 
# A:- 11111111111111111111111111111001
# A:- 11111111111111111111111111100100
# -----------------------------------------------
# --------> a>>>=2 <-------- 
# A:- 11111111111111111111111111111001
# A:- 11111111111111111111111111111110
# -----------------------------------------------
# 	--> ADD A:- 30 | B:- 60 || C:- 90
# 	--> SUB A:- 60 | B:- 20 || C:- 40
# 	--> MUL A:- 30 | B:- 60 || C:- 1800
# 	--> DIV A:- 30 | B:- 5 || C:- 6
# 	--> MOD A:- 30 | B:- 5 || C:- 0
# 	--> POW A:- 2 | B:- 12 || C:- 4096
# -----------------------------------------------
# 	--> AND A:- 1011 B:- 11 C:- 11
# 	--> OR A:- 1011 B:- 11 C:- 1011
# 	--> NAND A:- 1011 B:- 11 C:- 11111111111111111111111111111100
# 	--> NOR A:- 1011 B:- 11 C:- 11111111111111111111111111110100
# 	--> XOR A:- 1011 B:- 11 C:- 1000
# 	--> XNOR A:- 1011 B:- 11 C:- 11111111111111111111111111110111
# 	--> NOT A:- 1011 C:- 11111111111111111111111111110100
# 	--> NOT B:- 11 C:- 11111111111111111111111111111100
# -----------------------------------------------
# 	--> LOGICAL_AND A:- 1000 B:- 0 C:- 0
# 	--> LOGICAL_!AND A:- 1000 B:- 0 C:- 1
# 	--> LOGICAL_OR A:- 1000 B:- 0 C:- 1
# 	--> LOGICAL_!OR A:- 1000 B:- 0 C:- 0
# -----------------------------------------------
*/
