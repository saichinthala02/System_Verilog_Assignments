module top;
	int intA[100],intA1[200];
	int varr;
	bit exist_f;
	initial begin
		varr=1322;
		for(int i=0;i<200;i++)begin
			intA1[i]=$urandom_range(200,999);
		end
		foreach(intA[i]) intA[i]=$urandom_range(999,1999);

		$display("Array-1(intA):- %p",intA);
		$display("-------------------------------------------------------------------");
		$display("Array-2(intA1):- %p",intA1);
		$display("-------------------------------------------------------------------");
		$display("\t--> Checking Without membership Operator <--");
		foreach(intA1[i])begin
			if(varr==intA[i] || varr==intA1[i]) exist_f=1;
		end
		if(exist_f==1) $display("\tvarr=%0d is present in any one of the Array",varr);
		else $display("\tvarr=%0d is not present in any one of the Array",varr); 
		$display("-------------------------------------------------------------------");
		$display("\t--> Checking using Membership Operator <--");
		if(varr inside {intA,intA1}) exist_f=1;
		else exist_f =0;
		if(exist_f==1) $display("\tvarr=%0d is present in any one of the Array",varr);
		else $display("\tvarr=%0d is not present in any one of the Array",varr); 
		$display("-------------------------------------------------------------------");
	end
endmodule

/* Output:-
# Start time: 16:24:09 on Nov 03,2025
# Array-1(intA):- '{1016, 1935, 1879, 1876, 1460, 1132, 1817, 1831, 1659, 1172, 1489, 1885, 1976, 1113, 1209, 1477, 1387, 1322, 1466, 1834, 1454, 1202, 1364, 1305, 1877, 1299, 1504, 1800, 1862, 1723, 1121, 1047, 1160, 1679, 1457, 1723, 1499, 1841, 1366, 1622, 1441, 1651, 1843, 1800, 1477, 1366, 1059, 1637, 1042, 1700, 1694, 1712, 1744, 1676, 1887, 1419, 1134, 1267, 1194, 1841, 1378, 1271, 1937, 1971, 1225, 1241, 1631, 1034, 1044, 1070, 1221, 1733, 1345, 1763, 1450, 1230, 1111, 1950, 1729, 1098, 1214, 1565, 1420, 1082, 1901, 1012, 1239, 1581, 1779, 1201, 1405, 1930, 1725, 1778, 1223, 1790, 1980, 1309, 1263, 1657}
# -------------------------------------------------------------------
# Array-2(intA1):- '{512, 590, 942, 862, 846, 590, 922, 822, 591, 258, 658, 828, 855, 382, 573, 764, 502, 421, 611, 749, 555, 776, 493, 269, 493, 529, 517, 818, 480, 595, 446, 209, 961, 488, 968, 630, 764, 438, 296, 607, 301, 655, 544, 217, 698, 299, 412, 859, 450, 334, 542, 813, 626, 951, 407, 652, 497, 979, 687, 815, 730, 585, 301, 984, 862, 325, 442, 638, 963, 296, 509, 249, 955, 328, 415, 933, 252, 645, 770, 396, 959, 433, 210, 253, 326, 756, 422, 939, 624, 644, 291, 827, 695, 447, 819, 911, 680, 209, 978, 681, 364, 904, 855, 439, 717, 981, 372, 952, 497, 964, 589, 879, 387, 486, 777, 525, 470, 840, 765, 744, 364, 275, 720, 389, 756, 325, 979, 530, 713, 634, 958, 878, 412, 457, 700, 745, 520, 913, 814, 508, 454, 306, 848, 619, 791, 340, 358, 974, 432, 525, 582, 460, 925, 693, 638, 677, 359, 801, 257, 393, 245, 517, 215, 409, 237, 322, 600, 208, 510, 950, 316, 352, 409, 580, 885, 201, 351, 622, 952, 495, 987, 388, 510, 656, 298, 782, 801, 539, 311, 476, 463, 944, 883, 602, 914, 694, 884, 327, 751, 313}
# -------------------------------------------------------------------
# 	--> Checking Without membership Operator <--
# 	varr=1322 is present in any one of the Array
# -------------------------------------------------------------------
# 	--> Checking using Membership Operator <--
# 	varr=1322 is present in any one of the Array
# -------------------------------------------------------------------
*/
