//--> Q2. Using Streaming Operator,push data into Queue.
module top;
	typedef logic unsigned [3:0] nibble;
	byte byteQ[$];
	bit [127:0] data;
	nibble nibbleQ[$];
	integer seed;
	initial begin
		data=$random;
		$display("Data:- %0d",data);
		$display("Data:- %0b",data);
		$display("-----------------------------------------------------------------------------------------------------------");
		$display("--> Byte Queue <--");
		byteQ = {>>byte{data}};
		$display("Right Streaming Queue:- %p",byteQ);
		byteQ = {<<byte{data}};
		$display("Left Streaming Queue:- %p",byteQ);
		$display("-----------------------------------------------------------------------------------------------------------");
		$display("-----------------------------------------------------------------------------------------------------------");
		$display("--> Nibble Queue <--");
		nibbleQ = {>>nibble{data}};
		$display("Right Streaming Queue:- %p",nibbleQ);
		nibbleQ = {<<nibble{data}};
		$display("Left Streaming Queue:- %p",nibbleQ);
		$display("-----------------------------------------------------------------------------------------------------------");
	end
endmodule

/* Output:-
# Start time: 17:25:00 on Nov 03,2025
# Data:- 303379748
# Data:- 00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000101010011010100100100
# -----------------------------------------------------------------------------------------------------------
# --> Byte Queue <--
# Right Streaming Queue:- '{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 21, 53, 36}
# Left Streaming Queue:- '{36, 53, 21, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0}
# -----------------------------------------------------------------------------------------------------------
# -----------------------------------------------------------------------------------------------------------
# --> Nibble Queue <--
# Right Streaming Queue:- '{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 5, 3, 5, 2, 4}
# Left Streaming Queue:- '{4, 2, 5, 3, 5, 1, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0}
# -----------------------------------------------------------------------------------------------------------
================================================================================================================================
# Data:- 127
# Data:- 1111111
# -----------------------------------------------------------------------------------------------------------
# --> Byte Queue <--
# Right Streaming Queue:- '{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 127}
# Left Streaming Queue:- '{127, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0}
# -----------------------------------------------------------------------------------------------------------
# -----------------------------------------------------------------------------------------------------------
# --> Nibble Queue <--
# Right Streaming Queue:- '{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 15}
# Left Streaming Queue:- '{15, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0}
# -----------------------------------------------------------------------------------------------------------
*/
