//--> Q9. Diff b/w unary and Arthmetic Operators.
--> Unary Operators

Definition: Operators that act on a single operand (one variable or value).
Purpose: They perform operations like increment, decrement, negation, or logical NOT.
Examples:
	int a = 5;
	int b = -a;   // Unary minus: makes it negative → b = -5
	int c = +a;   // Unary plus: keeps it same → c = 5
	a++;          // Increment → a = 6
	a--;          // Decrement → a = 5
	
--> Arithmetic Operators
Definition: Operators that perform mathematical operations between two operands.
Purpose: Used for standard arithmetic calculations.
Examples:	
	int a = 10, b = 3;
	int sum = a + b;   // Addition → 13
	int diff = a - b;  // Subtraction → 7
	int prod = a * b;  // Multiplication → 30
	int div = a / b;   // Division → 3
	int mod = a % b;   // Modulus → 1


//--> Q10. Practical applications of unary operators
--> Loop control / Iteration
--> Address pointer updates
--> Signed arithmetic operations
--> Signal polarity inversion
--> Conditional control logic
--> Active-low signal generation
--> Bit masking / Bit inversion
--> Parity generation
--> Error detection / Bus integrity check
	
