//--> Q16. Multidimensional Array.
module top;
	reg [7:0][9:0] multi_arr[8][6:0];
	initial begin
		for(int i=0;i<8;i++)begin
			for(int j=0;j<7;j++)begin
				for(int k=0;k<8;k++)begin
					multi_arr[i][j][k]=$urandom_range(0,1023);
					$display("multi_arr[%0d][%0d][%0d]=%0d",i,j,k,multi_arr[i][j][k]);   
				end
			end
		end
		$display("The Array Elements:- %p",multi_arr);
	end
endmodule

/* Output:-
# Start time: 19:21:44 on Oct 31,2025
# The Array Elements:- '{'{'{68, 239, 783, 490, 613, 502, 742, 602}, '{435, 852, 547, 306, 337, 600, 967, 293}, '{407, 192, 398, 212, 526, 896, 320, 697}, '{969, 342, 395, 344, 394, 93, 745, 293}, '{773, 485, 800, 739, 517, 987, 381, 174}, '{980, 565, 598, 623, 436, 106, 314, 103}, '{814, 882, 582, 198, 950, 358, 38, 952}}, '{'{167, 741, 508, 169, 720, 876, 973, 325}, '{367, 943, 864, 516, 705, 618, 265, 256}, '{743, 267, 439, 559, 755, 411, 444, 904}, '{707, 510, 588, 254, 725, 266, 137, 951}, '{132, 410, 989, 980, 29, 343, 160, 883}, '{657, 693, 832, 731, 790, 466, 285, 630}, '{816, 901, 993, 498, 711, 839, 203, 457}}, '{'{936, 880, 410, 613, 1009, 719, 733, 109}, '{545, 633, 505, 287, 125, 630, 13, 373}, '{676, 1022, 709, 328, 70, 894, 1004, 431}, '{3, 552, 202, 638, 1012, 518, 873, 352}, '{33, 980, 737, 212, 582, 342, 690, 353}, '{426, 683, 893, 620, 701, 168, 907, 452}, '{0, 277, 928, 910, 389, 673, 190, 59}}, '{'{170, 493, 200, 896, 448, 513, 478, 757}, '{430, 30, 140, 427, 195, 860, 593, 852}, '{340, 1000, 790, 292, 405, 623, 234, 1013}, '{145, 711, 479, 44, 334, 394, 82, 1003}, '{200, 359, 436, 943, 883, 569, 294, 834}, '{712, 150, 828, 371, 295, 752, 582, 695}, '{193, 845, 636, 593, 280, 436, 1006, 886}}, '{'{39, 983, 690, 924, 81, 252, 564, 60}, '{361, 322, 975, 490, 719, 425, 503, 783}, '{522, 267, 923, 395, 423, 274, 531, 65}, '{422, 646, 272, 409, 976, 718, 17, 91}, '{480, 390, 480, 1022, 932, 918, 278, 400}, '{731, 300, 72, 797, 565, 437, 83, 943}, '{591, 424, 354, 286, 182, 884, 345, 805}}, '{'{356, 297, 922, 629, 406, 535, 51, 914}, '{848, 310, 710, 784, 819, 200, 674, 10}, '{700, 929, 696, 496, 139, 336, 248, 812}, '{813, 845, 596, 924, 646, 909, 919, 755}, '{985, 396, 832, 544, 347, 271, 736, 949}, '{257, 533, 139, 468, 942, 847, 257, 370}, '{329, 213, 157, 19, 251, 449, 595, 417}}, '{'{625, 906, 225, 765, 75, 414, 357, 274}, '{881, 193, 965, 32, 490, 619, 796, 892}, '{952, 421, 515, 440, 62, 107, 22, 583}, '{795, 869, 209, 668, 826, 229, 684, 156}, '{951, 714, 551, 402, 56, 836, 539, 211}, '{539, 696, 879, 724, 1000, 866, 481, 994}, '{395, 73, 617, 964, 363, 56, 536, 988}}, '{'{993, 871, 746, 155, 488, 777, 665, 921}, '{974, 1022, 985, 421, 752, 894, 2, 287}, '{86, 99, 486, 222, 806, 802, 315, 879}, '{884, 438, 3, 17, 632, 134, 499, 639}, '{27, 819, 513, 563, 305, 862, 327, 736}, '{354, 280, 31, 896, 244, 260, 731, 535}, '{762, 876, 977, 523, 717, 791, 477, 115}}}
----------------------------------------------------------------------------------------------------------------------------------------
# multi_arr[0][0][0]=952
# multi_arr[0][0][1]=38
# multi_arr[0][0][2]=358
# multi_arr[0][0][3]=950
# multi_arr[0][0][4]=198
# multi_arr[0][0][5]=582
# multi_arr[0][0][6]=882
# multi_arr[0][0][7]=814
# multi_arr[0][1][0]=103
# multi_arr[0][1][1]=314
# multi_arr[0][1][2]=106
# multi_arr[0][1][3]=436
# multi_arr[0][1][4]=623
# multi_arr[0][1][5]=598
# multi_arr[0][1][6]=565
# multi_arr[0][1][7]=980
# multi_arr[0][2][0]=174
# multi_arr[0][2][1]=381
# multi_arr[0][2][2]=987
# multi_arr[0][2][3]=517
# multi_arr[0][2][4]=739
# multi_arr[0][2][5]=800
# multi_arr[0][2][6]=485
# multi_arr[0][2][7]=773
# multi_arr[0][3][0]=293
# multi_arr[0][3][1]=745
# multi_arr[0][3][2]=93
# multi_arr[0][3][3]=394
# multi_arr[0][3][4]=344
# multi_arr[0][3][5]=395
# multi_arr[0][3][6]=342
# multi_arr[0][3][7]=969
# multi_arr[0][4][0]=697
# multi_arr[0][4][1]=320
# multi_arr[0][4][2]=896
# multi_arr[0][4][3]=526
# multi_arr[0][4][4]=212
# multi_arr[0][4][5]=398
# multi_arr[0][4][6]=192
# multi_arr[0][4][7]=407
# multi_arr[0][5][0]=293
# multi_arr[0][5][1]=967
# multi_arr[0][5][2]=600
# multi_arr[0][5][3]=337
# multi_arr[0][5][4]=306
# multi_arr[0][5][5]=547
# multi_arr[0][5][6]=852
# multi_arr[0][5][7]=435
# multi_arr[0][6][0]=602
# multi_arr[0][6][1]=742
# multi_arr[0][6][2]=502
# multi_arr[0][6][3]=613
# multi_arr[0][6][4]=490
# multi_arr[0][6][5]=783
# multi_arr[0][6][6]=239
# multi_arr[0][6][7]=68
# multi_arr[1][0][0]=457
# multi_arr[1][0][1]=203
# multi_arr[1][0][2]=839
# multi_arr[1][0][3]=711
# multi_arr[1][0][4]=498
# multi_arr[1][0][5]=993
# multi_arr[1][0][6]=901
# multi_arr[1][0][7]=816
# multi_arr[1][1][0]=630
# multi_arr[1][1][1]=285
# multi_arr[1][1][2]=466
# multi_arr[1][1][3]=790
# multi_arr[1][1][4]=731
# multi_arr[1][1][5]=832
# multi_arr[1][1][6]=693
# multi_arr[1][1][7]=657
# multi_arr[1][2][0]=883
# multi_arr[1][2][1]=160
# multi_arr[1][2][2]=343
# multi_arr[1][2][3]=29
# multi_arr[1][2][4]=980
# multi_arr[1][2][5]=989
# multi_arr[1][2][6]=410
# multi_arr[1][2][7]=132
# multi_arr[1][3][0]=951
# multi_arr[1][3][1]=137
# multi_arr[1][3][2]=266
# multi_arr[1][3][3]=725
# multi_arr[1][3][4]=254
# multi_arr[1][3][5]=588
# multi_arr[1][3][6]=510
# multi_arr[1][3][7]=707
# multi_arr[1][4][0]=904
# multi_arr[1][4][1]=444
# multi_arr[1][4][2]=411
# multi_arr[1][4][3]=755
# multi_arr[1][4][4]=559
# multi_arr[1][4][5]=439
# multi_arr[1][4][6]=267
# multi_arr[1][4][7]=743
# multi_arr[1][5][0]=256
# multi_arr[1][5][1]=265
# multi_arr[1][5][2]=618
# multi_arr[1][5][3]=705
# multi_arr[1][5][4]=516
# multi_arr[1][5][5]=864
# multi_arr[1][5][6]=943
# multi_arr[1][5][7]=367
# multi_arr[1][6][0]=325
# multi_arr[1][6][1]=973
# multi_arr[1][6][2]=876
# multi_arr[1][6][3]=720
# multi_arr[1][6][4]=169
# multi_arr[1][6][5]=508
# multi_arr[1][6][6]=741
# multi_arr[1][6][7]=167
# multi_arr[2][0][0]=59
# multi_arr[2][0][1]=190
# multi_arr[2][0][2]=673
# multi_arr[2][0][3]=389
# multi_arr[2][0][4]=910
# multi_arr[2][0][5]=928
# multi_arr[2][0][6]=277
# multi_arr[2][0][7]=0
# multi_arr[2][1][0]=452
# multi_arr[2][1][1]=907
# multi_arr[2][1][2]=168
# multi_arr[2][1][3]=701
# multi_arr[2][1][4]=620
# multi_arr[2][1][5]=893
# multi_arr[2][1][6]=683
# multi_arr[2][1][7]=426
# multi_arr[2][2][0]=353
# multi_arr[2][2][1]=690
# multi_arr[2][2][2]=342
# multi_arr[2][2][3]=582
# multi_arr[2][2][4]=212
# multi_arr[2][2][5]=737
# multi_arr[2][2][6]=980
# multi_arr[2][2][7]=33
# multi_arr[2][3][0]=352
# multi_arr[2][3][1]=873
# multi_arr[2][3][2]=518
# multi_arr[2][3][3]=1012
# multi_arr[2][3][4]=638
# multi_arr[2][3][5]=202
# multi_arr[2][3][6]=552
# multi_arr[2][3][7]=3
# multi_arr[2][4][0]=431
# multi_arr[2][4][1]=1004
# multi_arr[2][4][2]=894
# multi_arr[2][4][3]=70
# multi_arr[2][4][4]=328
# multi_arr[2][4][5]=709
# multi_arr[2][4][6]=1022
# multi_arr[2][4][7]=676
# multi_arr[2][5][0]=373
# multi_arr[2][5][1]=13
# multi_arr[2][5][2]=630
# multi_arr[2][5][3]=125
# multi_arr[2][5][4]=287
# multi_arr[2][5][5]=505
# multi_arr[2][5][6]=633
# multi_arr[2][5][7]=545
# multi_arr[2][6][0]=109
# multi_arr[2][6][1]=733
# multi_arr[2][6][2]=719
# multi_arr[2][6][3]=1009
# multi_arr[2][6][4]=613
# multi_arr[2][6][5]=410
# multi_arr[2][6][6]=880
# multi_arr[2][6][7]=936
# multi_arr[3][0][0]=886
# multi_arr[3][0][1]=1006
# multi_arr[3][0][2]=436
# multi_arr[3][0][3]=280
# multi_arr[3][0][4]=593
# multi_arr[3][0][5]=636
# multi_arr[3][0][6]=845
# multi_arr[3][0][7]=193
# multi_arr[3][1][0]=695
# multi_arr[3][1][1]=582
# multi_arr[3][1][2]=752
# multi_arr[3][1][3]=295
# multi_arr[3][1][4]=371
# multi_arr[3][1][5]=828
# multi_arr[3][1][6]=150
# multi_arr[3][1][7]=712
# multi_arr[3][2][0]=834
# multi_arr[3][2][1]=294
# multi_arr[3][2][2]=569
# multi_arr[3][2][3]=883
# multi_arr[3][2][4]=943
# multi_arr[3][2][5]=436
# multi_arr[3][2][6]=359
# multi_arr[3][2][7]=200
# multi_arr[3][3][0]=1003
# multi_arr[3][3][1]=82
# multi_arr[3][3][2]=394
# multi_arr[3][3][3]=334
# multi_arr[3][3][4]=44
# multi_arr[3][3][5]=479
# multi_arr[3][3][6]=711
# multi_arr[3][3][7]=145
# multi_arr[3][4][0]=1013
# multi_arr[3][4][1]=234
# multi_arr[3][4][2]=623
# multi_arr[3][4][3]=405
# multi_arr[3][4][4]=292
# multi_arr[3][4][5]=790
# multi_arr[3][4][6]=1000
# multi_arr[3][4][7]=340
# multi_arr[3][5][0]=852
# multi_arr[3][5][1]=593
# multi_arr[3][5][2]=860
# multi_arr[3][5][3]=195
# multi_arr[3][5][4]=427
# multi_arr[3][5][5]=140
# multi_arr[3][5][6]=30
# multi_arr[3][5][7]=430
# multi_arr[3][6][0]=757
# multi_arr[3][6][1]=478
# multi_arr[3][6][2]=513
# multi_arr[3][6][3]=448
# multi_arr[3][6][4]=896
# multi_arr[3][6][5]=200
# multi_arr[3][6][6]=493
# multi_arr[3][6][7]=170
# multi_arr[4][0][0]=805
# multi_arr[4][0][1]=345
# multi_arr[4][0][2]=884
# multi_arr[4][0][3]=182
# multi_arr[4][0][4]=286
# multi_arr[4][0][5]=354
# multi_arr[4][0][6]=424
# multi_arr[4][0][7]=591
# multi_arr[4][1][0]=943
# multi_arr[4][1][1]=83
# multi_arr[4][1][2]=437
# multi_arr[4][1][3]=565
# multi_arr[4][1][4]=797
# multi_arr[4][1][5]=72
# multi_arr[4][1][6]=300
# multi_arr[4][1][7]=731
# multi_arr[4][2][0]=400
# multi_arr[4][2][1]=278
# multi_arr[4][2][2]=918
# multi_arr[4][2][3]=932
# multi_arr[4][2][4]=1022
# multi_arr[4][2][5]=480
# multi_arr[4][2][6]=390
# multi_arr[4][2][7]=480
# multi_arr[4][3][0]=91
# multi_arr[4][3][1]=17
# multi_arr[4][3][2]=718
# multi_arr[4][3][3]=976
# multi_arr[4][3][4]=409
# multi_arr[4][3][5]=272
# multi_arr[4][3][6]=646
# multi_arr[4][3][7]=422
# multi_arr[4][4][0]=65
# multi_arr[4][4][1]=531
# multi_arr[4][4][2]=274
# multi_arr[4][4][3]=423
# multi_arr[4][4][4]=395
# multi_arr[4][4][5]=923
# multi_arr[4][4][6]=267
# multi_arr[4][4][7]=522
# multi_arr[4][5][0]=783
# multi_arr[4][5][1]=503
# multi_arr[4][5][2]=425
# multi_arr[4][5][3]=719
# multi_arr[4][5][4]=490
# multi_arr[4][5][5]=975
# multi_arr[4][5][6]=322
# multi_arr[4][5][7]=361
# multi_arr[4][6][0]=60
# multi_arr[4][6][1]=564
# multi_arr[4][6][2]=252
# multi_arr[4][6][3]=81
# multi_arr[4][6][4]=924
# multi_arr[4][6][5]=690
# multi_arr[4][6][6]=983
# multi_arr[4][6][7]=39
# multi_arr[5][0][0]=417
# multi_arr[5][0][1]=595
# multi_arr[5][0][2]=449
# multi_arr[5][0][3]=251
# multi_arr[5][0][4]=19
# multi_arr[5][0][5]=157
# multi_arr[5][0][6]=213
# multi_arr[5][0][7]=329
# multi_arr[5][1][0]=370
# multi_arr[5][1][1]=257
# multi_arr[5][1][2]=847
# multi_arr[5][1][3]=942
# multi_arr[5][1][4]=468
# multi_arr[5][1][5]=139
# multi_arr[5][1][6]=533
# multi_arr[5][1][7]=257
# multi_arr[5][2][0]=949
# multi_arr[5][2][1]=736
# multi_arr[5][2][2]=271
# multi_arr[5][2][3]=347
# multi_arr[5][2][4]=544
# multi_arr[5][2][5]=832
# multi_arr[5][2][6]=396
# multi_arr[5][2][7]=985
# multi_arr[5][3][0]=755
# multi_arr[5][3][1]=919
# multi_arr[5][3][2]=909
# multi_arr[5][3][3]=646
# multi_arr[5][3][4]=924
# multi_arr[5][3][5]=596
# multi_arr[5][3][6]=845
# multi_arr[5][3][7]=813
# multi_arr[5][4][0]=812
# multi_arr[5][4][1]=248
# multi_arr[5][4][2]=336
# multi_arr[5][4][3]=139
# multi_arr[5][4][4]=496
# multi_arr[5][4][5]=696
# multi_arr[5][4][6]=929
# multi_arr[5][4][7]=700
# multi_arr[5][5][0]=10
# multi_arr[5][5][1]=674
# multi_arr[5][5][2]=200
# multi_arr[5][5][3]=819
# multi_arr[5][5][4]=784
# multi_arr[5][5][5]=710
# multi_arr[5][5][6]=310
# multi_arr[5][5][7]=848
# multi_arr[5][6][0]=914
# multi_arr[5][6][1]=51
# multi_arr[5][6][2]=535
# multi_arr[5][6][3]=406
# multi_arr[5][6][4]=629
# multi_arr[5][6][5]=922
# multi_arr[5][6][6]=297
# multi_arr[5][6][7]=356
# multi_arr[6][0][0]=988
# multi_arr[6][0][1]=536
# multi_arr[6][0][2]=56
# multi_arr[6][0][3]=363
# multi_arr[6][0][4]=964
# multi_arr[6][0][5]=617
# multi_arr[6][0][6]=73
# multi_arr[6][0][7]=395
# multi_arr[6][1][0]=994
# multi_arr[6][1][1]=481
# multi_arr[6][1][2]=866
# multi_arr[6][1][3]=1000
# multi_arr[6][1][4]=724
# multi_arr[6][1][5]=879
# multi_arr[6][1][6]=696
# multi_arr[6][1][7]=539
# multi_arr[6][2][0]=211
# multi_arr[6][2][1]=539
# multi_arr[6][2][2]=836
# multi_arr[6][2][3]=56
# multi_arr[6][2][4]=402
# multi_arr[6][2][5]=551
# multi_arr[6][2][6]=714
# multi_arr[6][2][7]=951
# multi_arr[6][3][0]=156
# multi_arr[6][3][1]=684
# multi_arr[6][3][2]=229
# multi_arr[6][3][3]=826
# multi_arr[6][3][4]=668
# multi_arr[6][3][5]=209
# multi_arr[6][3][6]=869
# multi_arr[6][3][7]=795
# multi_arr[6][4][0]=583
# multi_arr[6][4][1]=22
# multi_arr[6][4][2]=107
# multi_arr[6][4][3]=62
# multi_arr[6][4][4]=440
# multi_arr[6][4][5]=515
# multi_arr[6][4][6]=421
# multi_arr[6][4][7]=952
# multi_arr[6][5][0]=892
# multi_arr[6][5][1]=796
# multi_arr[6][5][2]=619
# multi_arr[6][5][3]=490
# multi_arr[6][5][4]=32
# multi_arr[6][5][5]=965
# multi_arr[6][5][6]=193
# multi_arr[6][5][7]=881
# multi_arr[6][6][0]=274
# multi_arr[6][6][1]=357
# multi_arr[6][6][2]=414
# multi_arr[6][6][3]=75
# multi_arr[6][6][4]=765
# multi_arr[6][6][5]=225
# multi_arr[6][6][6]=906
# multi_arr[6][6][7]=625
# multi_arr[7][0][0]=115
# multi_arr[7][0][1]=477
# multi_arr[7][0][2]=791
# multi_arr[7][0][3]=717
# multi_arr[7][0][4]=523
# multi_arr[7][0][5]=977
# multi_arr[7][0][6]=876
# multi_arr[7][0][7]=762
# multi_arr[7][1][0]=535
# multi_arr[7][1][1]=731
# multi_arr[7][1][2]=260
# multi_arr[7][1][3]=244
# multi_arr[7][1][4]=896
# multi_arr[7][1][5]=31
# multi_arr[7][1][6]=280
# multi_arr[7][1][7]=354
# multi_arr[7][2][0]=736
# multi_arr[7][2][1]=327
# multi_arr[7][2][2]=862
# multi_arr[7][2][3]=305
# multi_arr[7][2][4]=563
# multi_arr[7][2][5]=513
# multi_arr[7][2][6]=819
# multi_arr[7][2][7]=27
# multi_arr[7][3][0]=639
# multi_arr[7][3][1]=499
# multi_arr[7][3][2]=134
# multi_arr[7][3][3]=632
# multi_arr[7][3][4]=17
# multi_arr[7][3][5]=3
# multi_arr[7][3][6]=438
# multi_arr[7][3][7]=884
# multi_arr[7][4][0]=879
# multi_arr[7][4][1]=315
# multi_arr[7][4][2]=802
# multi_arr[7][4][3]=806
# multi_arr[7][4][4]=222
# multi_arr[7][4][5]=486
# multi_arr[7][4][6]=99
# multi_arr[7][4][7]=86
# multi_arr[7][5][0]=287
# multi_arr[7][5][1]=2
# multi_arr[7][5][2]=894
# multi_arr[7][5][3]=752
# multi_arr[7][5][4]=421
# multi_arr[7][5][5]=985
# multi_arr[7][5][6]=1022
# multi_arr[7][5][7]=974
# multi_arr[7][6][0]=921
# multi_arr[7][6][1]=665
# multi_arr[7][6][2]=777
# multi_arr[7][6][3]=488
# multi_arr[7][6][4]=155
# multi_arr[7][6][5]=746
# multi_arr[7][6][6]=871
# multi_arr[7][6][7]=993
*/

/*
e. multi_arr[6] : how many bits does it represent.
	row 6 has: 7 columns,8 locations, 10 bit size 
	total bits:- 7*8*10 ==> 560 bits.

f. multi_arr[6][2] : how many bits does it represent.
	total bits:- 8*10 ==> 80 bits.

g. multi_arr[6][2][1] : how many bits does it represent.
	total bits:- 10 bits.

h. multi_arr[6][2][1][4] : how many bits does it represent.
	total bits:- 1 bit.
*/	
