module top;
	typedef int que[$];
	typedef que da[];
	typedef da arr[10];
    arr a;

	initial begin
		for(int i=0;i<10;i++)begin
          a[i]=new[5];
          for(int j=0;j<5;j++)begin
				repeat(3)begin
                  a[i][j].push_back($urandom_range(10,15));
				end
			end
		end
		$display("arr=%p",a);
	end
endmodule

/* Output:-
# arr='{'{'{11, 12, 12}, '{13, 12, 10}, '{14, 14, 12}, '{12, 12, 13}, '{14, 11, 15}},
	    '{'{13, 10, 14}, '{10, 15, 12}, '{14, 12, 11}, '{10, 10, 14}, '{13, 15, 10}}, 
		'{'{10, 12, 13}, '{15, 12, 12}, '{12, 12, 11}, '{13, 13, 12}, '{10, 15, 13}}, 
		'{'{13, 12, 12}, '{13, 11, 11}, '{12, 14, 14}, '{11, 14, 15}, '{10, 15, 10}}, 
		'{'{14, 12, 13}, '{15, 15, 11}, '{11, 12, 14}, '{13, 12, 13}, '{15, 13, 15}}, 
		'{'{14, 14, 11}, '{13, 11, 13}, '{10, 11, 15}, '{12, 14, 15}, '{12, 12, 14}}, 
		'{'{13, 11, 14}, '{15, 13, 12}, '{13, 10, 15}, '{14, 14, 11}, '{14, 10, 11}}, 
		'{'{12, 11, 10}, '{12, 10, 14}, '{11, 11, 11}, '{12, 14, 13}, '{11, 11, 12}}, 
		'{'{14, 15, 10}, '{11, 15, 14}, '{15, 14, 12}, '{12, 12, 13}, '{14, 10, 11}}, 
		'{'{11, 10, 13}, '{10, 12, 13}, '{14, 14, 12}, '{12, 14, 10}, '{12, 10, 12}}}
*/
