class eth_bad_pkt extends eth_pkt;
	static int count_bad;

	function new();
		count_bad++;
	endfunction
	
	function void print(string str="eth_bad_pkt");
		super.print(str);
		$display("Count_Bad:- %0d",count_bad);
	endfunction
endclass
