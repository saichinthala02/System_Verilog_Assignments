class eth_ext_pkt extends eth_pkt;
	
endclass
